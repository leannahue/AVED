library IEEE;
use IEEE.std_logic_1164.all;

--Additional standard or custom libraries go here
package canny_constants is
	--constant IMG_WIDTH	: natural := 480;
	--constant IMG_HEIGHT	: natural := 480;
	constant IMG_WIDTH	: natural := 5;
	constant IMG_HEIGHT	: natural := 5;

	constant MAG_WIDTH	: natural := 10;
end package canny_constants;

package body canny_constants is

end package body canny_constants;


